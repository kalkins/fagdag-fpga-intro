module top(
   input        clk,
   input        rst_n,
   output [7:0] led
);

   // TODO

endmodule
